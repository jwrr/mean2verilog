module tb;


parameter WID = 16;

reg           clk;
reg           rst;
reg [WID-1:0] in_000;
reg [WID-1:0] in_001;
reg [WID-1:0] in_002;
reg [WID-1:0] in_003;
reg [WID-1:0] in_004;
reg [WID-1:0] in_005;
reg [WID-1:0] in_006;
reg [WID-1:0] in_007;

reg test_done;

mean8 u_mean8(
    .clk     (clk),
    .rst     (rst),
    .in_000  (in_000),
    .in_001  (in_001),
    .in_002  (in_002),
    .in_003  (in_003),
    .in_004  (in_004),
    .in_005  (in_005),
    .in_006  (in_006),
    .in_007  (in_007)
);


// ============================================================================
// ============================================================================


initial
 begin
    $dumpfile("tb_mean.vcd");
    $dumpvars(0,tb);
 end


// ============================================================================
// ============================================================================


initial begin
    clk <= 0;
    #10;
    while (!test_done) begin
        #5 clk <= !clk;
    end
end


// ============================================================================
// ============================================================================


task clkn(input integer n);
begin
    repeat(n)
        @(posedge clk);
end
endtask


// ============================================================================
// ============================================================================


initial begin
  test_done <= 0;
  rst    <= 0;
  in_000 <= 10;
  in_001 <= 11;
  in_002 <= 12;
  in_003 <= 13;
  in_004 <= 14;
  in_005 <= 15;
  in_006 <= 16;
  in_007 <= 17;


  $display($time);
  clkn(10);
  rst <= 1;
  clkn(10);
  rst <= 0;
  clkn(10);
  
  repeat(100) begin
      in_000 <= in_000 + 1;
      in_001 <= in_001 + 1;
      in_002 <= in_002 + 1;
      in_003 <= in_003 + 1;
      in_004 <= in_004 + 1;
      in_005 <= in_005 + 1;
      in_006 <= in_006 + 1;
      in_007 <= in_007 + 1;
      clkn(1);
  end

  $display($time);
  $finish();
end



endmodule

